
module clockslow (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
