module counter_register(input [31:0] val);
integer [31:0] value;

value = val;
endmodule
